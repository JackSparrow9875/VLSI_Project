4-bit full adder implementation

.include TSMC_180nm.txt
.include NAND.sub
.include OR.sub
.include AND.sub
.include XOR.sub
.include NOT.sub
.include full_adder.sub
.include 4-bit_adder.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a0 a0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_a1 a1 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_a2 a2 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_a3 a3 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)

V_in_b0 b0 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_b1 b1 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_b2 b2 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_b3 b3 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)

V_in_m m gnd dc 0

X1 a0 a1 a2 a3 b0 b1 b2 b3 m sum0 sum1 sum2 sum3 carry node_x gnd four_bit_adder

.tran 1n 800n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(a0) v(a1)+2 v(a2)+4 v(a3)+6
hardcopy adder_subtractor_a_inp v(a0) v(a1)+2 v(a2)+4 v(a3)+6
plot v(b0) v(b1)+2 v(b2)+4 v(b3)+6
hardcopy adder_subtractor_b_inp v(b0) v(b1)+2 v(b2)+4 v(b3)+6
plot v(sum0) v(sum1)+2 v(sum2)+4 v(sum3)+6
hardcopy adder_subtractor_output v(sum0) v(sum1)+2 v(sum2)+4 v(sum3)+6
.end
.endc