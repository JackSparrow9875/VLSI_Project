4-bit full adder implementation

.include TSMC_180nm.txt
.include NAND.sub
.include OR.sub
.include AND.sub
.include XOR.sub
.include NOT.sub
.include XNOR.sub
.include 4-bit_comparator.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a0 a0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_a1 a1 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_a2 a2 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_a3 a3 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)

V_in_b0 b0 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_b1 b1 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_b2 b2 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_b3 b3 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)

X1 a0 a1 a2 a3 b0 b1 b2 b3 greater equal lesser node_x gnd fourbit_comparator

.tran 1n 800n

.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(a0) v(a1)+2 v(a2)+4 v(a3)+6
plot v(b0) v(b1)+2 v(b2)+4 v(b3)+6
plot v(greater) v(equal)+2 v(lesser)+4 
.end
.endc