full adder implementation

.include TSMC_180nm.txt
.include NAND.sub
.include OR.sub
.include AND.sub
.include XOR.sub
.include NOT.sub
.include full_adder.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a node_a gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b node_b gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)
V_in_c node_c gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)

X1 node_a node_b node_c sum carry node_x gnd full_adder

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = black
plot v(node_a) v(node_b)+2 v(node_c)+4 v(sum)+6 v(carry)+8
.end
.endc